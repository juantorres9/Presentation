library verilog;
use verilog.vl_types.all;
entity fiabilitetp1_vlg_vec_tst is
end fiabilitetp1_vlg_vec_tst;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


ENTITY fiabilitetp1 IS
GENERIC(
N: INTEGER:=3
);
PORT(
--ENTREES
  A: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);--6=Rin  543=SWITCH A ----210=SWITCH B
  B: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);--ASSIGNATION X3 SWITCH B
  Rin: IN STD_LOGIC;
iCLK_50: IN STD_LOGIC;
iCLK_50_2: IN STD_LOGIC;

oHEX0_D: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);--LEDS 7 segments
--SORTIES
S: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0);--- 210=MAX SOMME SUR N bits 
Rout:OUT STD_LOGIC
);
END fiabilitetp1;

ARCHITECTURE arch2 OF fiabilitetp1 IS 
SIGNAL TOTAL : STD_LOGIC_VECTOR(N DOWNTO 0);--SIGNAL QUI STOCK LE RESULTAT AVEC DEPASSEMENT EN BIT 3

--COMPONENT
COMPONENT AFFICHEUR IS
PORT (
SW: IN STD_LOGIC_VECTOR( 3 downto 0);-- SWITCH physique de 0000 � 1111
HEX: OUT STD_LOGIC_VECTOR( 6 DOWNTO 0) -- sorties physique vers les afficheurs
);
END COMPONENT;

BEGIN
PROCESS
VARIABLE RinS:   STD_LOGIC_VECTOR(0 DOWNTO 0);
BEGIN
WAIT UNTIL iCLK_50 ='1';
RinS(0):=Rin;
TOTAL <=STD_LOGIC_VECTOR(UNSIGNED('0'&A(N-1 DOWNTO 0))+UNSIGNED(B(N-1 DOWNTO 0))+UNSIGNED(RinS));
END PROCESS;
S(N-1 DOWNTO 0)<=TOTAL(N-1 DOWNTO 0);--Affichage LEDS =3210
Rout<=TOTAL(N);------Affichage LED MSB=3

instance1:afficheur PORT MAP(SW=> STD_LOGIC_VECTOR(TOTAL),HEX=>oHEX0_D);
END arch2;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


ENTITY dff8 IS
GENERIC(
N: INTEGER:=8
);
PORT(
--ENTREES
D: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
CLK: IN STD_LOGIC;
--SORTIES
Q: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
);
END dff8;

ARCHITECTURE arch1 OF dff8 IS 
BEGIN
PROCESS
BEGIN
WAIT UNTIL CLK'EVENT AND CLK= '1';
Q <=D;
END PROCESS;
END arch1;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


ENTITY additioneur IS
GENERIC(
N: INTEGER:=3
);
PORT(
--ENTREES
A: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
B: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
Rin: IN STD_LOGIC;
CLK: IN STD_LOGIC;
--SORTIES
S: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0);
Rout:OUT STD_LOGIC
);
END additioneur;

ARCHITECTURE arch2 OF additioneur IS 
SIGNAL TOTAL : STD_LOGIC_VECTOR(N DOWNTO 0);--SIGNAL QUI STOCKE LE RESULTAT AVEC DEPASSEMENT EN BIT 9
BEGIN
PROCESS
VARIABLE RinS:   STD_LOGIC_VECTOR(0 DOWNTO 0);
BEGIN
WAIT UNTIL CLK ='1';
RinS(0):=Rin;
TOTAL <=STD_LOGIC_VECTOR(UNSIGNED('0'&A)+UNSIGNED(B)+UNSIGNED(RinS));
END PROCESS;
S<=TOTAL(N-1 DOWNTO 0);
Rout<=TOTAL(N);
END arch2;

library verilog;
use verilog.vl_types.all;
entity dff8_vlg_vec_tst is
end dff8_vlg_vec_tst;

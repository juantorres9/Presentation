LIBRARY IEEE; 
USE ieee.std_logic_1164.ALL; 

ENTITY ALU IS 
PORT(
A: STD_LOGIC_VECTOR(2 DOWNTO 0) 
)
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


ENTITY basculemulti IS
GENERIC(
N: INTEGER :=4
);
PORT(
--ENTREES
A: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);--0010  =2
B: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);--1101  =13 OU -3
SEL:IN STD_LOGIC_VECTOR(1 DOWNTO 0);
--SORTIES
C: OUT STD_LOGIC_VECTOR(2*N-1 DOWNTO 0)--00000000
);
END basculemulti;


ARCHITECTURE arch3 OF basculemulti IS  
SIGNAL C1,C4: SIGNED(2*N-1 DOWNTO 0);
SIGNAL C2,C3: UNSIGNED(2*N-1 DOWNTO 0);
BEGIN

PROCESS(SEL,A,B)
BEGIN
C1<=SIGNED(A)*SIGNED(B);--OPERATION     2*-3=-6=1111 1010 le systeme remplis de 1 le reste de  Bits jusque a ZERO
C2<=UNSIGNED(A)*UNSIGNED(B);--OPERATION 2*13=26 0001 1010
C3<=UNSIGNED(A&"00")+"00000000";--2*4=8=1000
C4(4 DOWNTO 0)<=SIGNED('0'&A)+SIGNED(B);--OPERATION   2+(-3)=-1=0000 1111
END PROCESS;

C<= STD_LOGIC_VECTOR(C1) WHEN SEL="00" ELSE
STD_LOGIC_VECTOR(C2) WHEN SEL="01" ELSE
STD_LOGIC_VECTOR(C3) WHEN SEL="10" ELSE
STD_LOGIC_VECTOR(C4) WHEN SEL="11" ;

END arch3;

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY afficheur IS
PORT(

SW:  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);-- INPUT Switch 4 Bits pour selectioner nombre de 0 a 15 
HEX: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)--OUTPUT 7 LEDS qui vont representer le nombre binaire a 4 bits 
);
END afficheur;


ARCHITECTURE archi OF afficheur IS 
SIGNAL HEXS: STD_LOGIC_VECTOR(6 DOWNTO 0);
BEGIN 

PROCESS(SW)
BEGIN


IF(SW="0000")THEN --Nombre 0
HEXS<="1000000";
ELSIF(SW="0001")THEN--Nombre 1
HEXS<="1111001";
ELSIF(SW="0010")THEN--Nombre 2
HEXS<="0100100";
ELSIF(SW="0011")THEN--Nombre 3
HEXS<="0110000";
ELSIF(SW="0100")THEN--Nombre 4
HEXS<="0011001";
ELSIF(SW="0101")THEN--Nombre 5
HEXS<="0010010";
ELSIF(SW="0110")THEN--Nombre 6
HEXS<="0000010";
ELSIF(SW="0111")THEN--Nombre 7
HEXS<="1111000";
ELSIF(SW="1000")THEN--Nombre 8
HEXS<="0000000";
ELSIF(SW="1001")THEN--Nombre 9
HEXS<="0010000";
ELSIF(SW="1010")THEN--Nombre A
HEXS<="0001000";
ELSIF(SW="1010")THEN--Nombre B
HEXS<="0000011";
ELSIF(SW="1011")THEN--Nombre C
HEXS<="1000110";
ELSIF(SW="1100")THEN--Nombre C
HEXS<="1000110";
ELSIF(SW="1101")THEN--Nombre D
HEXS<="0100001";
ELSIF(SW="1110")THEN--Nombre E
HEXS<="0000110";
ELSIF(SW="1111")THEN--Nombre F
HEXS<="0001110";
ELSE--Nombre Error
HEXS<="1111110";
END IF;

END PROCESS;
HEX<=HEXS;
END archi;
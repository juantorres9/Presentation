LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


ENTITY additioneur2 IS
GENERIC(
N: INTEGER:=1;--Bits pour representer  l'Addition A5=(2*N-1)  et B + Rin 
R: INTEGER:=3 --Bits pour representer la somme de 3 2 1 0=0 à F
);
PORT(
--ENTREES
iSW: IN STD_LOGIC_VECTOR(2*N DOWNTO 0);--2=Rin  1=SWITCH A ----0=SWITCH B
iCLK_50: IN STD_LOGIC;
oHEX0_D: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);--LEDS 7 segments
--SORTIES
oLEDG:   OUT STD_LOGIC_VECTOR(R DOWNTO 0)---3=Rout  210=MAX SOMME SUR N bits 
--Rout:OUT STD_LOGIC
);
END additioneur2;

ARCHITECTURE arch2 OF additioneur2 IS 
SIGNAL TOTAL : STD_LOGIC_VECTOR(R DOWNTO 0);--SIGNAL QUI STOCKE LE RESULTAT AVEC DEPASSEMENT EN BIT 4

--COMPONENT
COMPONENT AFFICHEUR IS
PORT (
SW: IN STD_LOGIC_VECTOR( R downto 0);-- SWITCH physique de 0000 a 1111
HEX: OUT STD_LOGIC_VECTOR( 6 DOWNTO 0) -- sorties physique vers les afficheurs
);
END COMPONENT;

BEGIN
PROCESS
VARIABLE RinS:   STD_LOGIC_VECTOR(0 DOWNTO 0);


BEGIN
WAIT UNTIL iCLK_50 ='1';
RinS(0):=iSW(2*N);
TOTAL <=STD_LOGIC_VECTOR(UNSIGNED("000"&iSW(2*N-1 DOWNTO N))+UNSIGNED(iSW(N-1 DOWNTO 0))+UNSIGNED(RinS));
END PROCESS;


oLEDG(R DOWNTO 0)<=TOTAL(R DOWNTO 0);--Affichage LEDS =3210
instance1:afficheur PORT MAP(SW=> STD_LOGIC_VECTOR(TOTAL),HEX=>oHEX0_D);
END arch2;

library verilog;
use verilog.vl_types.all;
entity parite_vlg_vec_tst is
end parite_vlg_vec_tst;
